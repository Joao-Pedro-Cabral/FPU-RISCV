
package config_pkg;

  localparam integer Exponent = 8;
  localparam integer Fraction = 23;

endpackage
